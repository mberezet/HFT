`define NODES 4
/*1 less than width*/
`define WORD_WIDTH 31
`define PRED_WIDTH 6
`define WEIGHT_WIDTH 24
