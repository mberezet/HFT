`ifndef _CONST_VH_
`define _CONST_VH_

`define NODES 6
/*1 less than width*/
`define VERT_WIDTH 39
`define WEIGHT_WIDTH 31
`define PRED_WIDTH 6

`end