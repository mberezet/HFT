'define NODES 66

module FOREX(input logic clk,
				input logic signal,
				input logic 