`define NODES 66
