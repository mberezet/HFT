`define NODES 1
