`define NODES 4
