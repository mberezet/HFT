//Comparator

module comp(input logic clk,
				input logic signal,
				input logic 