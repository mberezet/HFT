module FOREX();

endmodule
